pll_2_inst : pll_2 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
